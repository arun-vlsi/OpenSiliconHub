// -----------------------------------------------------------------------------
// Module: lcg (Linear Congruential Generator)
// Author: MrAbhi19
// Description:
//   This module implements a Linear Congruential Generator (LCG),
//   a pseudo-random number generator defined by the recurrence:
//       X_{n+1} = (A * X_n + C) mod M
//
//   Each clock cycle produces the next pseudo-random number in the sequence.
//   The generator is initialized with a seed value.
//
// Parameters:
//   A - Multiplier constant (default = 214013)
//   C - Increment constant (default = 2531011)
//   M - Modulus constant (default = 2^31)
//
//   ► Microsoft C Runtime (MSVCRT) Variant:
//     - A = 214013
//     - C = 2531011
//     - M = 2^31
//     This is the widely used LCG configuration in Microsoft's C standard library.
//     Using these values replicates the pseudo-random sequence generated by
//     the MSVCRT `rand()` function.
//
// Ports:
//   clk   - Input clock signal. Advances the generator on each rising edge.
//   rst   - Asynchronous reset. Resets the generator state to the seed.
//   seed  - 32-bit input seed value used to initialize the generator.
//           Valid range: 1 to (2^32 - 1).
//   out   - 32-bit output representing the current pseudo-random number.
//
// Notes:
//   - The modulo operator (%) may not synthesize efficiently for non-power-of-2 M.
//     For hardware optimization, consider restricting M to powers of 2.
//   - This design is sequential and requires a clock for proper operation.
//   - The output sequence is deterministic given the same seed and parameters.
// -----------------------------------------------------------------------------

module lcg #(
  parameter A = 214013,   // Multiplier constant (MSVCRT default)
  parameter C = 2531011,  // Increment constant (MSVCRT default)
  parameter M = 2**31     // Modulus constant (MSVCRT default)
)(
  input        clk,        // Clock input
  input        rst,        // Asynchronous reset input
  input  [30:0] seed,      // Seed value (1 to 2^32 - 1)
  output reg [30:0] out    // Current pseudo-random output
);

  reg [30:0] inter;        // Internal state register

  // Sequential logic: update state and output on clock or reset
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      inter <= seed;        // Initialize state with seed
      out   <= seed % M;    // Ensure output is within modulus range
    end else begin
      inter <= (inter * A + C) % M; // Compute next state
      out   <= inter;               // Update output
    end
  end

endmodule
